module
  input a 
