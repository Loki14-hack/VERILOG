module
  input a 


  
