module
  input a 

  
