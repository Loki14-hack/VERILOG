  module d_ff (
    input  wire clk,
    input  wire d,
    output reg  

    
